----------------------------------------------------------------------------------------
-- This file is part of the VISCY project.
-- (C) 2007-2021 Gundolf Kiefer, Fachhochschule Augsburg, University of Applied Sciences
-- (C) 2018 Michael SchÃ¤ferling, Hochschule Augsburg, University of Applied Sciences
--
-- Description:
--   This is a testbench for the VISCY CPU - neither exhaustive nor complete
----------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity VISCY_CPU_TB is
end VISCY_CPU_TB;


architecture BEHAVIOR of VISCY_CPU_TB is

  -- Component Declaration for the Unit Under Test (UUT) ...
  component CPU
    port (
      clk:    in    std_logic;
      reset:  in    std_logic;
      adr:    out   std_logic_vector (15 downto 0);
      rdata:  in    std_logic_vector (15 downto 0);
      wdata:  out   std_logic_vector (15 downto 0);
      rd:     out   std_logic;
      wr:     out   std_logic;
      ready:  in    std_logic
    );
  end component;

  -- Signals ...
  signal clk:   std_logic := '0';
  signal reset: std_logic := '0';
  signal ready: std_logic := '0';

  signal adr:   std_logic_vector(15 downto 0);
  signal rdata: std_logic_vector(15 downto 0);
  signal wdata: std_logic_vector(15 downto 0);
  signal rd:    std_logic;
  signal wr:    std_logic;

  -- Parameters...
  constant clk_period: time := 10 ns;
  constant mem_delay: time := 25 ns;

  -- Memory content (generated by viscy2l) ...

 type t_memory is array (0 to 71) of std_logic_vector (15 downto 0);
	signal mem_content: t_memory := (
      16#0000# => "0100100000000000",  -- LDIH  r0, 0x00   ; => 00000000
      16#0001# => "0100000000000000",  -- LDIL  r0, 0x00   ; => 0000000000000000
      16#0002# => "0100100100000000",  -- LDIH  r1, 0x00   ; => 00000000
      16#0003# => "0100000100000000",  -- LDIL  r1, 0x00   ; => 0000000000000000
      16#0004# => "0100101100000000",  -- LDIH  r3, 0x00   ; => 00000000
      16#0005# => "0100001100000000",  -- LDIL  r3, 0x00   ; => 0000000000000000
      16#0006# => "0100110000000000",  -- LDIH  r4, 0x00   ; => 00000000
      16#0007# => "0100011100000000",  -- LDIL  r7, 0x00   ; => 0000000000000000
      16#0008# => "0100111100000000",  -- LDIH  r7, 0x00   ; => 00000000
      16#0009# => "0100101000000000",  -- LDIH  r2, 0x00   ; => 00000000
      16#000a# => "0100001000000000",  -- LDIL  r2, 0x00   ; => 0000000000000000
      16#000b# => "0011000000000000",  -- XOR   r0, r0, r0 ; Nur '0' in r0   // bitweise XOR Operation zwischen den Register r0 und r0, wodurch Wert von r0 den Wert 0
      16#000c# => "0100000000010011",  -- LDIL  r0, 787      ; 1. Wert in r0.  //lädt das Immediate-Low-Byte des Wertes 8 in das Register r0
      16#000d# => "0011000100100100",  -- XOR   r1, r1, r1
      16#000e# => "0100000111100011",  -- LDIL  r1, 739
      16#000f# => "0011011111111100",  -- XOR   r7, r7, r7
      16#0010# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0011# => "0011010010010000",  -- XOR   r4, r4, r4
      16#0012# => "0000001100000100",  -- ADD   r3, r0, r1 ; Addition: r3 = r0 + r1     => 1526       addiert die Werte in den Registern r0 und r1 und speichert Ergebnis in r3
      16#0013# => "0100010011110110",  -- LDIL  r4, 1526
      16#0014# => "0011011101110000",  -- XOR   r7, r3, r4
      16#0015# => "0010101001011100",  -- OR    r2, r2, r7
      16#0016# => "0011010010010000",  -- XOR   r4, r4, r4
      16#0017# => "0011011111111100",  -- XOR   r7, r7, r7
      16#0018# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0019# => "0000101100000100",  -- SUB   r3, r0, r1 ; Subtraktion: r3 = r0 - r1  => 48
      16#001a# => "0100010000110000",  -- LDIL  r4, 48
      16#001b# => "0011011101110000",  -- XOR   r7, r3, r4
      16#001c# => "0010101001011100",  -- OR    r2, r2, r7
      16#001d# => "0011010010010000",  -- XOR   r4, r4, r4
      16#001e# => "0011011111111100",  -- XOR   r7, r7, r7
      16#001f# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0020# => "0001001100000000",  -- SAL   r3, r0     ; Links-Shift:               => 1574        Linksverschiebung (Shift) des Werts in Register r0 und speichert das Ergebnis in r3
      16#0021# => "0100010000100110",  -- LDIL  r4, 1574
      16#0022# => "0011011101110000",  -- XOR   r7, r3, r4
      16#0023# => "0010101001011100",  -- OR    r2, r2, r7
      16#0024# => "0011010010010000",  -- XOR   r4, r4, r4
      16#0025# => "0011011111111100",  -- XOR   r7, r7, r7
      16#0026# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0027# => "0001101100000000",  -- SAR   r3, r0     ; Rechts-Shift:              => 393
      16#0028# => "0100010010001001",  -- LDIL  r4, 393
      16#0029# => "0011011101110000",  -- XOR   r7, r3, r4
      16#002a# => "0010101001011100",  -- OR    r2, r2, r7
      16#002b# => "0011001101101100",  -- XOR   r3, r3, r3
      16#002c# => "0011010010010000",  -- XOR   r4, r4, r4
      16#002d# => "0011011111111100",  -- XOR   r7, r7, r7
      16#002e# => "0010001100000100",  -- AND   r3, r0, r1 ; => 721
      16#002f# => "0100010011010001",  -- LDIL  r4, 721
      16#0030# => "0011011101110000",  -- XOR   r7, r3, r4
      16#0031# => "0010101001011100",  -- OR    r2, r2, r7
      16#0032# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0033# => "0011010010010000",  -- XOR   r4, r4, r4
      16#0034# => "0011011111111100",  -- XOR   r7, r7, r7
      16#0035# => "0010101100000100",  -- OR    r3, r0, r1 ; => 795
      16#0036# => "0100010000011011",  -- LDIL  r4, 795
      16#0037# => "0011011101110000",  -- XOR   r7, r3, r4
      16#0038# => "0010101001011100",  -- OR    r2, r2, r7
      16#0039# => "0011001101101100",  -- XOR   r3, r3, r3
      16#003a# => "0011010010010000",  -- XOR   r4, r4, r4
      16#003b# => "0011011111111100",  -- XOR   r7, r7, r7
      16#003c# => "0011001100000100",  -- XOR   r3, r0, r1 ; => 64
      16#003d# => "0100010001000000",  -- LDIL  r4, 64
      16#003e# => "0011011101110000",  -- XOR   r7, r3, r4
      16#003f# => "0010101001011100",  -- OR    r2, r2, r7
      16#0040# => "0011001101101100",  -- XOR   r3, r3, r3
      16#0041# => "0011010010010000",  -- XOR   r4, r4, r4
      16#0042# => "0011011111111100",  -- XOR   r7, r7, r7
      16#0043# => "0011101100000000",  -- NOT   r3, r0     ; =>  476         bitweise Negation (NOT-Operation) des Werts in Register
      16#0044# => "0100010011011100",  -- LDIL  r4, 476
      16#0045# => "0011011101110000",  -- XOR   r7, r3, r4
      16#0046# => "0010101001011100",  -- OR    r2, r2, r7
      16#0047# => "1000100000000000",  -- HALT
      others => "UUUUUUUUUUUUUUUU"
    );


	for ALL: CPU use entity WORK.CPU(RTL);

BEGIN

  -- Instantiate the Unit Under Test (UUT)
  UUT: CPU port map (
      clk => clk,
      reset => reset,
      adr => adr,
      rdata => rdata,
      wdata => wdata,
      rd => rd,
      wr => wr,
      ready => ready
    );

  -- Process to simulate the memory behavior ...
  memory: process
  begin
    ready <= '0';
    wait on rd, wr;
    if rd = '1' then
      wait for mem_delay;
      if is_x (adr) then
        rdata <= (others => 'X');
      else
        rdata <= mem_content (to_integer (unsigned (adr)));
      end if;
      ready <= '1';
      wait until rd = '0';
      rdata <= (others => 'X');
      wait for mem_delay;
      ready <= '0';
    elsif wr = '1' then
      wait for mem_delay;
      if not is_x(adr) then
        mem_content (to_integer (unsigned (adr))) <= wdata;
      end if;
      ready <= '1';
      wait until wr = '0';
      wait for mem_delay;
      ready <= '0';
    end if;
  end process;


  -- Main testbench process ...
  testbench: process
    
    procedure run_cycle is
    begin
      clk <= '0';
      wait for clk_period / 2;
      clk <= '1';
      wait for clk_period / 2;
    end procedure;

    variable n: integer;
    
    variable memread: std_logic_vector(15 downto 0);
    
  begin

    -- HIER: SINNVOLLES HAUPTPROGRAMM EINFÃœGEN

    reset <= '1';
    run_cycle;
    reset <= '0';

    
    -- run cycle in while-loop until rd != '1' for 10 iterations (means that CPU stoppped => halt)
    n := 0;
    while n < 10 loop
		run_cycle;

		if rd = '0' then
			n := n + 1;
		else
			n := 0;
		end if;
	end loop;
        
    wait; -- wait forever (stop simulation)
  end process;

end;
